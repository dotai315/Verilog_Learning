module hello_world();
  initial begin
    $display("Hello World!");
  end
endmodule