module initial_example();

reg clk, reset, enable, data;

initial begin
  clk     = 0;
  reset   = 0;
  enable  = 0;
  data    = 0;
end

endmodule